`timescale 1ns/1ns
module IFstage
	(
		input clk,
		input rst,
		input br_taken,
		input [31:0]br_addr,
		output reg [31:0] PC_out,
		output [31:0] Instruction
	);
	
reg [31:0] PC_in = 32'd0;

wire[31 : 0]instMem[118 : 0];
assign instMem[0] = 32'b000000_00000_00000_00000_00000000000;//--NOP
//assign instMem[4] = 32'b100000_00000_00001_00000_11000001010;//-- Addi	r1	,r0	,1546
//assign instMem[8] = 32'b000011_00000_00001_00011_00000000000;//-- sub	r3	,r0	,r1 
//assign instMem[12] = 32'b000101_00010_00011_00100_00000000000;//-- And	r4	,r2	,r3	
//assign instMem[16] = 32'b100001_00011_00101_00011_01000110100;//-- Subi	r5	,r3	,6708   
//assign instMem[20] = 32'b000110_00011_00100_00101_00000000000;//-- or	r5	,r3	,r4
assign instMem[1] = 32'b100000_00000_00001_00000_11000001010;//-- Addi r1 ,r0 ,1546
assign instMem[2] = 32'b000000_00000_00000_00000_00000000000;//--NOP
assign instMem[3] = 32'b000000_00000_00000_00000_00000000000;//--NOP
assign instMem[4] = 32'b000000_00000_00000_00000_00000000000;//--NOP
assign instMem[5] = 32'b000001_00000_00001_00010_00000000000;//-- Add r2 ,r0 ,r1
assign instMem[6] = 32'b000011_00000_00001_00011_00000000000;//-- sub r3 ,r0 ,r1
assign instMem[7] = 32'b000000_00000_00000_00000_00000000000;//--NOP
assign instMem[8] = 32'b000000_00000_00000_00000_00000000000;//--NOP
assign instMem[9] = 32'b000000_00000_00000_00000_00000000000;//--NOP
assign instMem[10] = 32'b000101_00010_00011_00100_00000000000;//-- And r4 ,r2 ,r3
assign instMem[11] = 32'b100001_00011_00101_00011_01000110100;//-- Subi r5 ,r3 ,6708
assign instMem[12] = 32'b000000_00000_00000_00000_00000000000;//--NOP
assign instMem[13] = 32'b000000_00000_00000_00000_00000000000;//--NOP
assign instMem[14] = 32'b000110_00011_00100_00101_00000000000;//-- or r5 ,r3 ,r4
assign instMem[15] = 32'b000000_00000_00000_00000_00000000000;//--NOP
assign instMem[16] = 32'b000000_00000_00000_00000_00000000000;//--NOP
assign instMem[17] = 32'b000000_00000_00000_00000_00000000000;//--NOP
assign instMem[18] = 32'b000111_00101_00000_00110_00000000000;//-- nor r6 ,r5 ,r0
assign instMem[19] = 32'b000111_00100_00000_01011_00000000000;//-- nor r11 ,r4 ,r0
assign instMem[20] = 32'b000011_00101_00101_00101_00000000000;//-- sub r5 ,r5 ,r5
assign instMem[21] = 32'b100000_00000_00001_00000_10000000000;//-- Addi r1 ,r0 ,1024
assign instMem[22] = 32'b000000_00000_00000_00000_00000000000;//--NOP
assign instMem[23] = 32'b000000_00000_00000_00000_00000000000;//--NOP
assign instMem[24] = 32'b000000_00000_00000_00000_00000000000;//--NOP
assign instMem[25] = 32'b100101_00001_00010_00000_00000000000;//-- st r2 ,r1 ,0
assign instMem[26] = 32'b100100_00001_00101_00000_00000000000;//-- ld r5 ,r1 ,0
assign instMem[27] = 32'b000000_00000_00000_00000_00000000000;//--NOP
assign instMem[28] = 32'b000000_00000_00000_00000_00000000000;//--NOP
assign instMem[29] = 32'b101000_00101_00000_00000_00000000001;//-- Bez r5 ,1
assign instMem[30] = 32'b001000_00101_00001_00111_00000000000;//-- xor r7 ,r5 ,r1
assign instMem[31] = 32'b001000_00101_00001_00000_00000000000;//-- xor r0 ,r5 ,r1
assign instMem[32] = 32'b001001_00011_01011_00111_00000000000;//-- sla r7 ,r3 ,r11
assign instMem[33] = 32'b001010_00011_01011_01000_00000000000;//-- sll r8 ,r3 ,r11
assign instMem[34] = 32'b001011_00011_00100_01001_00000000000;//-- sra r9 ,r3 ,r4
assign instMem[35] = 32'b001100_00011_00100_01010_00000000000;//-- srl r10 ,r3 ,r4
assign instMem[36] = 32'b100101_00001_00011_00000_00000000100;//-- st r3 ,r1 ,4
assign instMem[37] = 32'b100101_00001_00100_00000_00000001000;//-- st r4 ,r1 ,8
assign instMem[38] = 32'b100101_00001_00101_00000_00000001100;//-- st r5 ,r1 ,12
assign instMem[39] = 32'b100101_00001_00110_00000_00000010000;//-- st r6 ,r1 ,16
assign instMem[40] = 32'b100100_00001_01011_00000_00000000100;//-- ld r11 ,r1 ,4
assign instMem[41] = 32'b100101_00001_00111_00000_00000010100;//-- st r7 ,r1 ,20
assign instMem[42] = 32'b100101_00001_01000_00000_00000011000;//-- st r8 ,r1 ,24
assign instMem[43] = 32'b100101_00001_01001_00000_00000011100;//-- st r9 ,r1 ,28
assign instMem[44] = 32'b100101_00001_01010_00000_00000100000;//-- st r10 ,r1 ,32
assign instMem[45] = 32'b100101_00001_01011_00000_00000100100;//-- st r11 ,r1 ,36
assign instMem[46] = 32'b100000_00000_00001_00000_00000000011;//-- Addi r1 ,r0 ,3
assign instMem[47] = 32'b100000_00000_00100_00000_10000000000;//-- Addi r4 ,r0 ,1024
assign instMem[48] = 32'b100000_00000_00010_00000_00000000000;//-- Addi r2 ,r0 ,0
assign instMem[49] = 32'b100000_00000_00011_00000_00000000001;//-- Addi r3 ,r0 ,1
assign instMem[50] = 32'b100000_00000_01001_00000_00000000010;//-- Addi r9 ,r0 ,2 	///////////
assign instMem[51] = 32'b000000_00000_00000_00000_00000000000;//--NOP
assign instMem[52] = 32'b000000_00000_00000_00000_00000000000;//--NOP
assign instMem[53] = 32'b000000_00000_00000_00000_00000000000;//--NOP
assign instMem[54] = 32'b001010_00011_01001_01000_00000000000;//-- sll r8 ,r3 ,r9
assign instMem[55] = 32'b000000_00000_00000_00000_00000000000;//--NOP
assign instMem[56] = 32'b000000_00000_00000_00000_00000000000;//--NOP
assign instMem[57] = 32'b000000_00000_00000_00000_00000000000;//--NOP
assign instMem[58] = 32'b000001_00100_01000_01000_00000000000;//-- Add r8 ,r4 ,r8
assign instMem[59] = 32'b000000_00000_00000_00000_00000000000;//--NOP
assign instMem[60] = 32'b000000_00000_00000_00000_00000000000;//--NOP
assign instMem[61] = 32'b000000_00000_00000_00000_00000000000;//--NOP
assign instMem[62] = 32'b100100_01000_00101_00000_00000000000;//-- ld r5 ,r8 ,0
assign instMem[63] = 32'b100100_01000_00110_11111_11111111100;//-- ld r6 ,r8 ,-4
assign instMem[64] = 32'b000000_00000_00000_00000_00000000000;//--NOP
assign instMem[65] = 32'b000000_00000_00000_00000_00000000000;//--NOP
assign instMem[66] = 32'b000000_00000_00000_00000_00000000000;//--NOP
assign instMem[67] = 32'b000011_00101_00110_01001_00000000000;//-- sub r9 ,r5 ,r6
assign instMem[68] = 32'b100000_00000_01010_10000_00000000000;//-- Addi r10 ,r0 ,0x8000
assign instMem[69] =  32'b100000_00000_01011_00000_00000010000;//-- Addi r11 ,r0 ,16
assign instMem[70] = 32'b000000_00000_00000_00000_00000000000;//--NOP
assign instMem[71] = 32'b000000_00000_00000_00000_00000000000;//--NOP
assign instMem[72] = 32'b000000_00000_00000_00000_00000000000;//--NOP
assign instMem[73] =  32'b001010_01010_01011_01010_00000000000;//-- sll r10 ,r1 ,r11
assign instMem[74] = 32'b000000_00000_00000_00000_00000000000;//--NOP
assign instMem[75] = 32'b000000_00000_00000_00000_00000000000;//--NOP
assign instMem[76] = 32'b000000_00000_00000_00000_00000000000;//--NOP
assign instMem[77] =  32'b000101_01001_01010_01001_00000000000;//-- And r9 ,r9 ,r10
assign instMem[78] = 32'b000000_00000_00000_00000_00000000000;//--NOP
assign instMem[79] = 32'b000000_00000_00000_00000_00000000000;//--NOP
assign instMem[80] = 32'b000000_00000_00000_00000_00000000000;//--NOP
assign instMem[81] =  32'b101000_01001_00000_00000_00000000010;//-- Bez r9 ,2
assign instMem[82] = 32'b000000_00000_00000_00000_00000000000;//--NOP
assign instMem[83] = 32'b000000_00000_00000_00000_00000000000;//--NOP
assign instMem[84] =  32'b100101_01000_00101_11111_11111111100;//-- st r5 ,r8 ,-4
assign instMem[85] =  32'b100101_01000_00110_00000_00000000000;//-- st r6 ,r8 ,0
assign instMem[86] =  32'b100000_00011_00011_00000_00000000001;//-- Addi r3 ,r3 ,1
assign instMem[87] = 32'b000000_00000_00000_00000_00000000000;//--NOP
assign instMem[88] = 32'b000000_00000_00000_00000_00000000000;//--NOP
assign instMem[89] = 32'b000000_00000_00000_00000_00000000000;//--NOP
assign instMem[90] = 32'b101001_00001_00011_11111_11111011000;//-- BNE r1 ,r3 ,-41		/////////////////////
assign instMem[91] = 32'b000000_00000_00000_00000_00000000000;//--NOP
assign instMem[92] = 32'b000000_00000_00000_00000_00000000000;//--NOP
assign instMem[93] =  32'b100000_00010_00010_00000_00000000001;//-- Addi r2 ,r2 ,1
assign instMem[94] = 32'b000000_00000_00000_00000_00000000000;//--NOP
assign instMem[95] = 32'b000000_00000_00000_00000_00000000000;//--NOP
assign instMem[96] = 32'b000000_00000_00000_00000_00000000000;//--NOP
assign instMem[97] =  32'b101001_00001_00010_11111_11111101110;//-- BNE r1 ,r2 ,-18
assign instMem[98] = 32'b000000_00000_00000_00000_00000000000;//--NOP
assign instMem[99] = 32'b000000_00000_00000_00000_00000000000;//--NOP
assign instMem[100] =  32'b100000_00000_00001_00000_10000000000;//-- Addi r1 ,r0 ,1024
assign instMem[101] = 32'b000000_00000_00000_00000_00000000000;//--NOP
assign instMem[102] = 32'b000000_00000_00000_00000_00000000000;//--NOP
assign instMem[103] = 32'b000000_00000_00000_00000_00000000000;//--NOP
assign instMem[104] =  32'b100100_00001_00010_00000_00000000000;//-- ld ,r2 ,r1 ,0
assign instMem[105] =  32'b100100_00001_00011_00000_00000000100;//-- ld ,r3 ,r1 ,4
assign instMem[106] =  32'b100100_00001_00100_00000_00000001000;//-- ld ,r4 ,r1 ,8
assign instMem[107] =  32'b100100_00001_00100_00000_01000001000;//-- ld ,r4 ,r1 ,520
assign instMem[108] =  32'b100100_00001_00100_00000_10000001000;//-- ld ,r4 ,r1 ,1023
assign instMem[109] =  32'b100100_00001_00101_00000_00000001100;//-- ld ,r5 ,r1 ,12
assign instMem[110] =  32'b100100_00001_00110_00000_00000010000;//-- ld ,r6 ,r1 ,16
assign instMem[111] =  32'b100100_00001_00111_00000_00000010100;//-- ld ,r7 ,r1 ,20
assign instMem[112] =  32'b100100_00001_01000_00000_00000011000;//-- ld ,r8 ,r1 ,24
assign instMem[113] =  32'b100100_00001_01001_00000_00000011100;//-- ld ,r9 ,r1 ,28
assign instMem[114] =  32'b100100_00001_01010_00000_00000100000;//-- ld ,r10,r1 ,32
assign instMem[115] =  32'b100100_00001_01011_00000_00000100100;//-- ld ,r11,r1 ,36
assign instMem[116] =  32'b101010_00000_00000_11111_11111111111;//-- JMP -1
assign instMem[117] = 32'b000000_00000_00000_00000_00000000000;//--NOP
assign instMem[118] = 32'b000000_00000_00000_00000_00000000000;//--NOP
assign instMem[118] = 32'b000000_00000_00000_00000_00000000000;//--NOP

	always@(posedge clk, posedge rst)begin
		if(rst)begin
			PC_out <= 32'd0;
		end
		else begin
			PC_out <= (br_taken)? br_addr : PC_out + 3'b100;
		end
	end
//assign PC_out = PC_in;
assign Instruction =(PC_out==0)? 32'b000000_00000_00000_00000_00000000000 : instMem[PC_out>>2];
endmodule
